32382
2014-04-17T00:00:00.000Z
-1609166.9529525214
884149.5805921489
-6939032.899708027
-2994.949034019323
6642.288367747897
1539.3798925236513
0.0
0.0
0.0
-1609166.9529525214
884149.5805921489
-6939032.899708027
-2994.949034019323
6642.288367747897
1539.3798925236513
0.0
0.0
0.0
2014-04-17T00:02:00.000Z
-1954811.120250542
1671353.49792403
-6701344.703493115
-2764.5992637523195
6476.936425853835
2421.597086097745
0.0
0.0
0.0
-1954811.120250542
1671353.49792403
-6701344.703493115
-2764.5992637523195
6476.936425853835
2421.597086097745
0.0
0.0
0.0
2014-04-17T00:04:00.000Z
-2270263.20692304
2432695.8418588648
-6360027.042530282
-2491.4898632706218
6211.438772165329
3266.357046284816
0.0
0.0
0.0
-2270263.20692304
2432695.8418588648
-6360027.042530282
-2491.4898632706218
6211.438772165329
3266.357046284816
0.0
0.0
0.0
2014-04-17T00:06:00.000Z
-2550642.8063140805
3156403.914758551
-5920356.180563221
-2179.821315312042
5849.883038741044
4060.645945769987
0.0
0.0
0.0
-2550642.8063140805
3156403.914758551
-5920356.180563221
-2179.821315312042
5849.883038741044
4060.645945769987
0.0
0.0
0.0
2014-04-17T00:08:00.000Z
-2791607.6092872648
3831282.439313085
-5389121.206097548
-1834.3834760586888
5397.822890102854
4792.217000659596
0.0
0.0
0.0
-2791607.6092872648
3831282.439313085
-5389121.206097548
-1834.3834760586888
5397.822890102854
4792.217000659596
0.0
0.0
0.0
2014-04-17T00:10:00.000Z
-2989423.4403111152
4446889.011933219
-4774529.118725438
-1460.4870731344008
4862.203579640577
5449.780587972664
0.0
0.0
0.0
-2989423.4403111152
4446889.011933219
-4774529.118725438
-1460.4870731344008
4862.203579640577
5449.780587972664
0.0
0.0
0.0
2014-04-17T00:12:00.000Z
-3141018.331830436
4993690.134582363
-4086071.6572899367
-1063.88118355755
4251.250605205363
6023.170174100957
0.0
0.0
0.0
-3141018.331830436
4993690.134582363
-4086071.6572899367
-1063.88118355755
4251.250605205363
6023.170174100957
0.0
0.0
0.0
2014-04-17T00:14:00.000Z
-3244029.7593986536
5463206.7413079515
-3334382.0608157134
-650.6678600638929
3574.348480446796
6503.496363678423
0.0
0.0
0.0
-3244029.7593986536
5463206.7413079515
-3334382.0608157134
-650.6678600638929
3574.348480446796
6503.496363678423
0.0
0.0
0.0
2014-04-17T00:16:00.000Z
-3296846.0125285205
5848152.21624123
-2531078.8342514886
-227.21205091534048
2841.9069618692233
6883.292330334122
0.0
0.0
0.0
-3296846.0125285205
5848152.21624123
-2531078.8342514886
-227.21205091534048
2841.9069618692233
6883.292330334122
0.0
0.0
0.0
2014-04-17T00:18:00.000Z
-3298627.539255819
6142538.64548673
-1688583.0783169332
199.95568406283104
2065.1998661076095
7156.622196171459
0.0
0.0
0.0
-3298627.539255819
6142538.64548673
-1688583.0783169332
199.95568406283104
2065.1998661076095
7156.622196171459
0.0
0.0
0.0
2014-04-17T00:20:00.000Z
-3249320.887217287
6341770.070666913
-819929.6868059845
624.2374812085583
1256.196882935002
7319.175044120566
0.0
0.0
0.0
-3249320.887217287
6341770.070666913
-819929.6868059845
624.2374812085583
1256.196882935002
7319.175044120566
0.0
0.0
0.0
2014-04-17T00:22:00.000Z
-3149665.4318655683
6442723.820845015
61429.59120577178
1039.0686310152614
427.3864429932369
7368.3455990790935
0.0
0.0
0.0
-3149665.4318655683
6442723.820845015
61429.59120577178
1039.0686310152614
427.3864429932369
7368.3455990790935
0.0
0.0
0.0
2014-04-17T00:24:00.000Z
-3001178.775025184
6443792.640810648
941835.5755367713
1438.018135796763
-408.41700817607693
7303.270068461865
0.0
0.0
0.0
-3001178.775025184
6443792.640810648
941835.5755367713
1438.018135796763
-408.41700817607693
7303.270068461865
0.0
0.0
0.0
2014-04-17T00:26:00.000Z
-2806134.933976055
6344911.979416495
1807630.6751045585
1814.887251499584
-1238.2672498481754
7124.84555158098
0.0
0.0
0.0
-2806134.933976055
6344911.979416495
1807630.6751045585
1814.887251499584
-1238.2672498481754
7124.84555158098
0.0
0.0
0.0
2014-04-17T00:28:00.000Z
-2567534.9592151637
6147573.015389634
2645371.325140711
2163.807847470577
-2049.2856926286436
6835.733266265953
0.0
0.0
0.0
-2567534.9592151637
6147573.015389634
2645371.325140711
2163.807847470577
-2049.2856926286436
6835.733266265953
0.0
0.0
0.0
2014-04-17T00:30:00.000Z
-2289057.276383859
5854793.102868265
3442036.787032396
2479.3331257128925
-2828.861807624027
6440.313415906151
0.0
0.0
0.0
-2289057.276383859
5854793.102868265
3442036.787032396
2479.3331257128925
-2828.861807624027
6440.313415906151
0.0
0.0
0.0
2014-04-17T00:32:00.000Z
-1975003.013519354
5471072.842757137
4185228.7696556565
2756.5225370112216
-3564.846799583327
5944.625222861342
0.0
0.0
0.0
-1975003.013519354
5471072.842757137
4185228.7696556565
2756.5225370112216
-3564.846799583327
5944.625222861342
0.0
0.0
0.0
2014-04-17T00:34:00.000Z
-1630232.9212800302
5002336.520350191
4863372.476064656
2991.0251581876255
-4245.7508273241465
5356.287454733238
0.0
0.0
0.0
-1630232.9212800302
5002336.520350191
4863372.476064656
2991.0251581876255
-4245.7508273241465
5356.287454733238
0.0
0.0
0.0
2014-04-17T00:36:00.000Z
-1260089.746609538
4455834.426525801
5465892.992779903
3179.146351526594
-4860.920773620349
4684.376330805737
0.0
0.0
0.0
-1260089.746609538
4455834.426525801
5465892.992779903
3179.146351526594
-4860.920773620349
4684.376330805737
0.0
0.0
0.0
2014-04-17T00:38:00.000Z
-870316.2085917068
3840032.7114031897
5983381.434725277
3317.908007201663
-5400.7098541674
3939.2890676252546
0.0
0.0
0.0
-870316.2085917068
3840032.7114031897
5983381.434725277
3317.908007201663
-5400.7098541674
3939.2890676252546
0.0
0.0
0.0
2014-04-17T00:40:00.000Z
-466967.66859719134
3164489.3107281066
6407751.984751619
3405.1025925353806
-5856.640154056166
3132.591223515113
0.0
0.0
0.0
-466967.66859719134
3164489.3107281066
6407751.984751619
3405.1025925353806
-5856.640154056166
3132.591223515113
0.0
0.0
0.0
2014-04-17T00:42:00.000Z
-56316.01836094301
2439699.663079076
6732363.05161466
3439.326168772231
-6221.533710515044
2276.8308003996394
0.0
0.0
0.0
-56316.01836094301
2439699.663079076
6732363.05161466
3439.326168772231
-6221.533710515044
2276.8308003996394
0.0
0.0
0.0
2014-04-17T00:44:00.000Z
355248.0614222145
1676933.9251837872
6952123.288090614
3420.0030243924593
-6489.629815711242
1385.3427015722618
0.0
0.0
0.0
355248.0614222145
1676933.9251837872
6952123.288090614
3420.0030243924593
-6489.629815711242
1385.3427015722618
0.0
0.0
0.0
2014-04-17T00:46:00.000Z
761314.9452437625
888064.854744805
7063582.860988488
3347.4019117520756
-6656.6888392667415
472.0425902578698
0.0
0.0
0.0
761314.9452437625
888064.854744805
7063582.860988488
3347.4019117520756
-6656.6888392667415
472.0425902578698
0.0
0.0
0.0
2014-04-17T00:48:00.000Z
1155557.2164489066
85377.77113271353
7064980.258690558
3222.628848635106
-6720.054588085578
-448.79756617183205
0.0
0.0
0.0
1155557.2164489066
85377.77113271353
7064980.258690558
3222.628848635106
-6720.054588085578
-448.79756617183205
0.0
0.0
0.0
2014-04-17T00:50:00.000Z
1531828.6517555383
-718621.1350742949
6956271.3632712085
3047.611165904621
-6678.699246478118
-1362.7751722542937
0.0
0.0
0.0
1531828.6517555383
-718621.1350742949
6956271.3632712085
3047.611165904621
-6678.699246478118
-1362.7751722542937
0.0
0.0
0.0
2014-04-17T00:52:00.000Z
1884263.0376826813
-1511402.0542499092
6739141.270353685
2825.072387735521
-6533.2515681597815
-2255.588299450706
0.0
0.0
0.0
1884263.0376826813
-1511402.0542499092
6739141.270353685
2825.072387735521
-6533.2515681597815
-2255.588299450706
0.0
0.0
0.0
2014-04-17T00:54:00.000Z
2207364.902969369
-2280608.6280364348
6416968.632058925
2558.484970285597
-6285.978759281274
-3113.263480190739
0.0
0.0
0.0
2207364.902969369
-2280608.6280364348
6416968.632058925
2558.484970285597
-6285.978759281274
-3113.263480190739
0.0
0.0
0.0
2014-04-17T00:56:00.000Z
2496095.9639869807
-3014252.131952914
5994772.92036521
2252.0152784094416
-5940.750949208865
-3922.378820135952
0.0
0.0
0.0
2496095.9639869807
-3014252.131952914
5994772.92036521
2252.0152784094416
-5940.750949208865
-3922.378820135952
0.0
0.0
0.0
2014-04-17T00:58:00.000Z
2745957.663973738
-3700903.6322771087
5479144.358575585
1910.4605821742414
-5502.988083685403
-4670.283246512555
0.0
0.0
0.0
2745957.663973738
-3700903.6322771087
5479144.358575585
1910.4605821742414
-5502.988083685403
-4670.283246512555
0.0
0.0
0.0
2014-04-17T01:00:00.000Z
2953058.8703624825
-4329870.8099655295
4878130.421393991
1539.168300091534
-4979.563255978147
-5345.294178409154
0.0
0.0
0.0
2953058.8703624825
-4329870.8099655295
4878130.421393991
1539.168300091534
-4979.563255978147
-5345.294178409154
0.0
0.0
0.0
2014-04-17T01:02:00.000Z
3114176.5420908337
-4891365.047190205
4201108.944227332
1143.9504659277577
-4378.691869887032
-5936.882230348606
0.0
0.0
0.0
3114176.5420908337
-4891365.047190205
4201108.944227332
1143.9504659277577
-4378.691869887032
-5936.882230348606
0.0
0.0
0.0
2014-04-17T01:04:00.000Z
3226810.0702532665
-5376660.449729171
3458647.138747547
730.9929054986966
-3709.8061967144913
-6435.8447205489065
0.0
0.0
0.0
3226810.0702532665
-5376660.449729171
3458647.138747547
730.9929054986966
-3709.8061967144913
-6435.8447205489065
0.0
0.0
0.0
2014-04-17T01:06:00.000Z
3289216.145469745
-5778225.255005796
2662325.507790568
306.7527889526412
-2983.394030836846
-6834.4435161821275
0.0
0.0
0.0
3289216.145469745
-5778225.255005796
2662325.507790568
306.7527889526412
-2983.394030836846
-6834.4435161821275
0.0
0.0
0.0
2014-04-17T01:08:00.000Z
3300434.766023565
-6089836.567540648
1824557.7263749545
-122.14290225351806
-2210.8321904227864
-7126.522398417459
0.0
0.0
0.0
3300434.766023565
-6089836.567540648
1824557.7263749545
-122.14290225351806
-2210.8321904227864
-7126.522398417459
0.0
0.0
0.0
2014-04-17T01:10:00.000Z
3260308.165271913
-6306685.18291203
958397.3744538378
-549.0031230022514
-1404.2068513741963
-7307.611010368801
0.0
0.0
0.0
3260308.165271913
-6306685.18291203
958397.3744538378
-549.0031230022514
-1404.2068513741963
-7307.611010368801
0.0
0.0
0.0
2014-04-17T01:12:00.000Z
3169477.413627911
-6425440.389497561
77328.8129057379
-967.1790331907963
-576.1162466006626
-7374.980479773329
0.0
0.0
0.0
3169477.413627911
-6425440.389497561
77328.8129057379
-967.1790331907963
-576.1162466006626
-7374.980479773329
0.0
0.0
0.0
2014-04-17T01:14:00.000Z
3029371.225476068
-6444299.224181216
-804942.899944883
-1370.167857221495
260.52811130892593
-7327.680387979028
0.0
0.0
0.0
3029371.225476068
-6444299.224181216
-804942.899944883
-1370.167857221495
260.52811130892593
-7327.680387979028
0.0
0.0
0.0
2014-04-17T01:16:00.000Z
2842186.729925904
-6363020.95189073
-1674706.7179038287
-1751.7160892386917
1092.705012827147
-7166.5577958467675
0.0
0.0
0.0
2842186.729925904
-6363020.95189073
-1674706.7179038287
-1751.7160892386917
1092.705012827147
-7166.5577958467675
0.0
0.0
0.0
2014-04-17T01:18:00.000Z
2610849.4446395454
-6182918.77357688
-2518459.0545859397
-2105.91483104554
1907.4880581191453
-6894.226861415893
0.0
0.0
0.0
2610849.4446395454
-6182918.77357688
-2518459.0545859397
-2105.91483104554
1907.4880581191453
-6894.226861415893
0.0
0.0
0.0
2014-04-17T01:20:00.000Z
2338966.6985885156
-5906836.539515313
-3323112.3847602997
-2427.290129416755
2692.2457524952497
-6515.021586891521
0.0
0.0
0.0
2338966.6985885156
-5906836.539515313
-3323112.3847602997
-2427.290129416755
2692.2457524952497
-6515.021586891521
0.0
0.0
0.0
2014-04-17T01:22:00.000Z
2030774.0213725474
-5539110.202619877
-4076201.0879087313
-2710.8892407639128
3434.8391893689004
-6034.931375623326
0.0
0.0
0.0
2030774.0213725474
-5539110.202619877
-4076201.0879087313
-2710.8892407639128
3434.8391893689004
-6034.931375623326
0.0
0.0
0.0
2014-04-17T01:24:00.000Z
1691064.6506250924
-5085488.968218447
-4766069.95559149
-2952.352269071706
4123.805161991458
-5461.492245167832
0.0
0.0
0.0
1691064.6506250924
-5085488.968218447
-4766069.95559149
-2952.352269071706
4123.805161991458
-5461.492245167832
0.0
0.0
0.0
2014-04-17T01:26:00.000Z
1325114.9641282056
-4553044.336431694
-5382051.556679956
-3147.9766069626544
4748.528847210775
-4803.665685802795
0.0
0.0
0.0
1325114.9641282056
-4553044.336431694
-5382051.556679956
-3147.9766069626544
4748.528847210775
-4803.665685802795
0.0
0.0
0.0
2014-04-17T01:28:00.000Z
938604.395679429
-3950065.330638674
-5914636.026991669
-3294.7755888086012
5299.409661413226
-4071.703033554219
0.0
0.0
0.0
938604.395679429
-3950065.330638674
-5914636.026991669
-3294.7755888086012
5299.409661413226
-4071.703033554219
0.0
0.0
0.0
2014-04-17T01:30:00.000Z
537525.0467187378
-3285921.7062551575
-6355608.619140934
-3390.517452726533
5767.9983501218485
-3276.9768493892702
0.0
0.0
0.0
537525.0467187378
-3285921.7062551575
-6355608.619140934
-3390.517452726533
5767.9983501218485
-3276.9768493892702
0.0
0.0
0.0
2014-04-17T01:32:00.000Z
128089.52479493678
-2570918.7980425917
-6698173.34703057
-3433.756778791624
6147.121325225072
-2431.804803474277
0.0
0.0
0.0
128089.52479493678
-2570918.7980425917
-6698173.34703057
-3433.756778791624
6147.121325225072
-2431.804803474277
0.0
0.0
0.0
2014-04-17T01:34:00.000Z
-283364.0212653265
-1816142.347520153
-6937064.001442938
-3423.858787136975
6430.993714181212
-1549.2640721834389
0.0
0.0
0.0
-283364.0212653265
-1816142.347520153
-6937064.001442938
-3423.858787136975
6430.993714181212
-1549.2640721834389
0.0
0.0
0.0
2014-04-17T01:36:00.000Z
-690469.949220154
-1033282.9687588578
-7068614.049573737
-3361.002176206275
6615.2952210116655
-642.9868345036481
0.0
0.0
0.0
-690469.949220154
-1033282.9687588578
-7068614.049573737
-3361.002176206275
6615.2952210116655
-642.9868345036481
0.0
0.0
0.0
2014-04-17T01:38:00.000Z
-1086932.159503665
-234457.23611906113
-7090810.625960102
-3246.174599426576
6697.231627065223
273.046048500138
0.0
0.0
0.0
-1086932.159503665
-234457.23611906113
-7090810.625960102
-3246.174599426576
6697.231627065223
273.046048500138
0.0
0.0
0.0
2014-04-17T01:40:00.000Z
-1466621.21181961
567976.5001218071
-7003333.570591863
-3081.1609538543426
6675.583084619873
1184.7155036731242
0.0
0.0
0.0
-1466621.21181961
567976.5001218071
-7003333.570591863
-3081.1609538543426
6675.583084619873
1184.7155036731242
0.0
0.0
0.0
2014-04-17T01:42:00.000Z
-1823667.1329948474
1361609.0057590194
-6807549.304464371
-2868.5107474522097
6550.711071973562
2077.9782782251727
0.0
0.0
0.0
-1823667.1329948474
1361609.0057590194
-6807549.304464371
-2868.5107474522097
6550.711071973562
2077.9782782251727
0.0
0.0
0.0
2014-04-17T01:44:00.000Z
-2152548.348889297
2134168.4539485043
-6506489.237855464
-2611.4993292700037
6324.551364307843
2939.076594100184
0.0
0.0
0.0
-2152548.348889297
2134168.4539485043
-6506489.237855464
-2611.4993292700037
6324.551364307843
2939.076594100184
0.0
0.0
0.0
DONE